module mux_4to1_2bitdata(
	output [1-0] out,
	input [1-0] in3,
	input [1-0] in2,
	input [1-0] in1,
	input [1-0] in0,
	);