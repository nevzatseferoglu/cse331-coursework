library verilog;
use verilog.vl_types.all;
entity Mips32_testbench is
end Mips32_testbench;
