
`define DELAY 20
module alu_32bit_testbench();

wire [31:0] r;
wire co;
wire z;

reg [2:0] aluOp;
reg [31:0] a;
reg [31:0] b;

alu_32bit test_alu (
	.r(r),
	.co(co),
	.z(z),
	
	.aluOp(aluOp),
	.a(a),
	.b(b)
	);

initial begin
	aluOp = 3'b000;
	a = 32'b 0000_0000_0000_0000_0000_0000_0000_0001;
	b = 32'b 0000_0000_0000_0000_0000_0000_0000_0001;
	#`DELAY;
	
	aluOp = 3'b000;
	a = 32'b 1000_0000_0000_0000_0000_0000_0000_0001;
	b = 32'b 0000_0000_0000_0000_0000_0000_0000_0000;
	#`DELAY;
	
	aluOp = 3'b001;
	a = 32'b 1000_0000_0000_0000_0000_0000_0000_0001;
	b = 32'b 0000_0000_0000_0000_0000_0000_0000_0000;
	#`DELAY;
	
	aluOp = 3'b001;
	a = 32'b 1111_0000_1111_0000_1111_0000_1111_0001;
	b = 32'b 0000_1111_0000_1111_0000_1111_0000_0000;
	#`DELAY;
	
	aluOp = 3'b010;
	a = 32'b 1111_1111_1111_1111_1111_1111_1111_1111;
	b = 32'b 1111_1111_1111_1111_1111_1111_1111_1111;
	#`DELAY;
	
	aluOp = 3'b110;
	a = 32'b 1111_1111_1111_1111_1111_1111_1111_1111;
	b = 32'b 1111_1111_1111_1111_1111_1111_1111_1111;
	#`DELAY;
	
	aluOp = 3'b110;
	a = 32'b 1111_1111_1111_1111_1111_1111_1111_1111;
	b = 32'b 0111_1111_1111_1111_1111_1111_1111_1111;
	#`DELAY;
	
	aluOp = 3'b011;
	a = 32'b 0000_0000_0000_0000_0000_0000_0000_0001;
	b = 32'b 0000_0000_0000_0000_0000_0000_0000_0001;
	#`DELAY;
	
	aluOp = 3'b011;
	a = 32'b 0101_1010_0000_0000_0000_0000_0000_0001;
	b = 32'b 1010_0101_0000_0000_0000_0000_0000_0000;
	#`DELAY;
	
end
 
 
initial begin
	$monitor("aluOp = %3b, a = %32b, b = %32b, result = %32b, co = %1b, z = %1b", aluOp, a, b, r, co, z);
end
 
endmodule




