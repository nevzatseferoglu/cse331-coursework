library verilog;
use verilog.vl_types.all;
entity Mips32 is
    port(
        clk             : in     vl_logic
    );
end Mips32;
