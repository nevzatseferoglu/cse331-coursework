module increment_by1_18bit (

);



endmodule
